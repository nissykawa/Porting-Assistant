* Created by KLayout

* cell Op8_22_rev2
* pin Bias
* pin In-
* pin In+
* pin Vdd
* pin Out
* pin Vss
.SUBCKT Op8_22_rev2 1 8 12 13 16 25
* net 1 Bias
* net 8 In-
* net 12 In+
* net 13 Vdd
* net 16 Out
* net 25 Vss
* device instance $1 m90 *1 35.5,41.5 NMOS
M$1 4 1 25 25 NMOS L=5U W=10U AS=15P AD=15P PS=21U PD=21U
* device instance $3 m90 *1 30.5,56 NMOS
M$3 11 1 4 25 NMOS L=2U W=20U AS=30P AD=30P PS=36U PD=36U
* device instance $5 m90 *1 96.5,61 NMOS
M$5 21 1 7 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $10 r0 *1 110.5,61 NMOS
M$10 10 1 3 25 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $15 r0 *1 142,42 NMOS
M$15 14 1 25 25 NMOS L=5U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $16 m90 *1 46,56 NMOS
M$16 1 1 6 25 NMOS L=2U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $17 m90 *1 95.5,41.5 NMOS
M$17 7 1 25 25 NMOS L=5U W=10U AS=15P AD=15P PS=21U PD=21U
* device instance $19 r0 *1 109.5,41.5 NMOS
M$19 3 1 25 25 NMOS L=5U W=10U AS=15P AD=15P PS=21U PD=21U
* device instance $21 r0 *1 59,41.5 NMOS
M$21 2 1 25 25 NMOS L=5U W=5U AS=10P AD=10P PS=14U PD=14U
* device instance $22 m90 *1 47.5,41.5 NMOS
M$22 6 1 25 25 NMOS L=5U W=5U AS=10P AD=10P PS=14U PD=14U
* device instance $23 r0 *1 55.5,56 NMOS
M$23 9 1 2 25 NMOS L=2U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $24 m0 *1 49.5,155.5 NMOS
M$24 11 8 24 25 NMOS L=3U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $28 r180 *1 37.5,155.5 NMOS
M$28 11 12 22 25 NMOS L=3U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $32 r0 *1 177,47 NMOS
M$32 16 10 25 25 NMOS L=1U W=96U AS=112P AD=112P PS=126U PD=126U
* device instance $38 m90 *1 167,49 NMOS
M$38 5 5 25 25 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $43 m90 *1 167,78 NMOS
M$43 15 15 5 25 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $48 m90 *1 165.5,111.5 NMOS
M$48 18 15 10 25 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $53 r0 *1 151.5,191.5 PMOS
M$53 15 9 13 13 PMOS L=5U W=16U AS=24P AD=24P PS=30U PD=30U
* device instance $55 m90 *1 99.5,185.5 PMOS
M$55 24 21 13 13 PMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $60 r0 *1 113,185.5 PMOS
M$60 22 21 13 13 PMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $65 m90 *1 90,152.5 PMOS
M$65 21 21 24 13 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $69 r0 *1 99.5,152.5 PMOS
M$69 18 21 22 13 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $73 r0 *1 52,188 PMOS
M$73 20 9 13 13 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $75 m90 *1 41,188 PMOS
M$75 23 9 13 13 PMOS L=5U W=15U AS=30P AD=30P PS=34U PD=34U
* device instance $76 r0 *1 190,165.5 PMOS
M$76 16 18 13 13 PMOS L=1U W=300U AS=420P AD=420P PS=434U PD=434U
* device instance $78 m90 *1 179,165.5 PMOS
M$78 19 19 13 13 PMOS L=1U W=300U AS=360P AD=360P PS=372U PD=372U
* device instance $83 m0 *1 31,123 PMOS
M$83 20 9 17 13 PMOS L=2U W=40U AS=60P AD=60P PS=66U PD=66U
* device instance $85 r180 *1 22,123 PMOS
M$85 23 9 9 13 PMOS L=2U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $86 m90 *1 143.5,98.5 PMOS
M$86 10 14 18 13 PMOS L=1U W=300U AS=330P AD=330P PS=352U PD=352U
* device instance $96 m90 *1 154.5,149 PMOS
M$96 14 14 19 13 PMOS L=1U W=300U AS=330P AD=330P PS=352U PD=352U
* device instance $106 m90 *1 70.5,104.5 PMOS
M$106 3 12 17 17 PMOS L=3U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $111 r0 *1 81.5,104.5 PMOS
M$111 7 8 17 17 PMOS L=3U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $119 r0 *1 7.5,179.5 HRES
R$119 1 13 800000 HRES
* device instance $124 r0 *1 289.25,49 CAP
C$124 16 10 1.4892e-12 CAP
* device instance $126 m0 *1 289.25,181 CAP
C$126 16 18 1.4892e-12 CAP
.ENDS Op8_22_rev2
