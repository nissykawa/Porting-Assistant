* Created by KLayout

* cell Op8_16_rev1
* pin Voutput
* pin Ibias1
* pin Vdd
* pin In+
* pin In-
* pin Vss
.SUBCKT Op8_16_rev1 7 8 10 15 16 17
* net 7 Voutput
* net 8 Ibias1
* net 10 Vdd
* net 15 In+
* net 16 In-
* net 17 Vss
* device instance $1 r0 *1 224.75,40.2 CAP
C$1 7 4 1.0366e-12 CAP
* device instance $5 r0 *1 55.5,100.5 NMOS
M$5 9 15 11 17 NMOS L=2U W=40U AS=80P AD=80P PS=84U PD=84U
* device instance $6 m90 *1 67.4,100.5 NMOS
M$6 12 16 11 17 NMOS L=2U W=40U AS=80P AD=80P PS=84U PD=84U
* device instance $7 m90 *1 17.1,18.1 NMOS
M$7 3 1 17 17 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $8 r0 *1 28,18.1 NMOS
M$8 2 1 17 17 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $9 r0 *1 113.5,23 NMOS
M$9 4 6 17 17 NMOS L=3U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $10 m90 *1 105,23 NMOS
M$10 6 6 17 17 NMOS L=3U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $11 r0 *1 64.7,36 NMOS
M$11 11 1 2 17 NMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $15 m90 *1 57.2,35.9 NMOS
M$15 1 1 3 17 NMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $19 r0 *1 126.3,19.35 NMOS
M$19 7 4 17 17 NMOS L=1U W=25U AS=37.5P AD=37.5P PS=43.5U PD=43.5U
* device instance $21 r0 *1 140.5,127.1 PMOS
M$21 7 8 10 10 PMOS L=5U W=90U AS=120P AD=120P PS=128U PD=128U
* device instance $24 r0 *1 121,127.1 PMOS
M$24 9 8 10 10 PMOS L=5U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $25 r0 *1 24,127 PMOS
M$25 14 8 10 10 PMOS L=5U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $26 m90 *1 13.1,127 PMOS
M$26 13 8 10 10 PMOS L=5U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $27 r0 *1 97.7,127.1 PMOS
M$27 12 8 10 10 PMOS L=5U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $28 r0 *1 22.6,82.9 PMOS
M$28 1 8 14 10 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $32 r0 *1 121.4,84.7 PMOS
M$32 4 8 9 10 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $36 r0 *1 87.5,84 PMOS
M$36 6 8 12 10 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $40 m90 *1 15,82.9 PMOS
M$40 8 8 13 10 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $44 r0 *1 -1,42 HRES
R$44 8 17 175000 HRES
.ENDS Op8_16_rev1
