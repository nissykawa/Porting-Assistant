* Created by KLayout

* cell Op8_22_rev2
* pin Bias
* pin In-
* pin In+
* pin Vdd
* pin Out
* pin Vss
.SUBCKT Op8_22_rev2 1 8 13 14 18 26
* net 1 Bias
* net 8 In-
* net 13 In+
* net 14 Vdd
* net 18 Out
* net 26 Vss
* device instance $1 m90 *1 35.5,41.5 NMOS
M$1 4 1 26 26 NMOS L=5U W=10U AS=15P AD=15P PS=21U PD=21U
* device instance $3 m90 *1 30.5,56 NMOS
M$3 12 1 4 26 NMOS L=2U W=20U AS=30P AD=30P PS=36U PD=36U
* device instance $5 r0 *1 142,42 NMOS
M$5 15 1 26 26 NMOS L=5U W=6U AS=15P AD=15P PS=17U PD=17U
* device instance $6 m90 *1 46,56 NMOS
M$6 1 1 6 26 NMOS L=2U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $7 r0 *1 109.5,41.5 NMOS
M$7 3 1 26 26 NMOS L=5U W=10U AS=15P AD=15P PS=21U PD=21U
* device instance $9 m90 *1 95.5,41.5 NMOS
M$9 7 1 26 26 NMOS L=5U W=10U AS=15P AD=15P PS=21U PD=21U
* device instance $11 r0 *1 59,41.5 NMOS
M$11 2 1 26 26 NMOS L=5U W=5U AS=10P AD=10P PS=14U PD=14U
* device instance $12 m90 *1 47.5,41.5 NMOS
M$12 6 1 26 26 NMOS L=5U W=5U AS=10P AD=10P PS=14U PD=14U
* device instance $13 r0 *1 55.5,56 NMOS
M$13 9 1 2 26 NMOS L=2U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $14 m90 *1 96.5,61 NMOS
M$14 10 1 7 26 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $19 r0 *1 110.5,61 NMOS
M$19 11 1 3 26 NMOS L=2U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $24 m0 *1 49.5,155.5 NMOS
M$24 12 8 25 26 NMOS L=3U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $28 r180 *1 37.5,155.5 NMOS
M$28 12 13 23 26 NMOS L=3U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $32 m90 *1 167,49 NMOS
M$32 5 5 26 26 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $37 m90 *1 167,78 NMOS
M$37 16 16 5 26 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $42 m90 *1 165.5,111.5 NMOS
M$42 20 16 11 26 NMOS L=1U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $47 r0 *1 177,47 NMOS
M$47 18 11 26 26 NMOS L=1U W=96U AS=112P AD=112P PS=126U PD=126U
* device instance $53 m90 *1 99.5,185.5 PMOS
M$53 25 10 14 14 PMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $58 r0 *1 113,185.5 PMOS
M$58 23 10 14 14 PMOS L=5U W=100U AS=120P AD=120P PS=132U PD=132U
* device instance $63 m90 *1 90,152.5 PMOS
M$63 10 10 25 14 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $67 r0 *1 99.5,152.5 PMOS
M$67 20 10 23 14 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $71 r0 *1 52,188 PMOS
M$71 22 9 14 14 PMOS L=5U W=30U AS=45P AD=45P PS=51U PD=51U
* device instance $73 m90 *1 41,188 PMOS
M$73 24 9 14 14 PMOS L=5U W=15U AS=30P AD=30P PS=34U PD=34U
* device instance $74 m90 *1 143.5,98.5 PMOS
M$74 11 15 20 14 PMOS L=1U W=300U AS=330P AD=330P PS=352U PD=352U
* device instance $84 m90 *1 154.5,149 PMOS
M$84 15 15 21 14 PMOS L=1U W=300U AS=330P AD=330P PS=352U PD=352U
* device instance $94 r0 *1 151.5,191.5 PMOS
M$94 16 9 14 14 PMOS L=5U W=16U AS=24P AD=24P PS=30U PD=30U
* device instance $96 r0 *1 190,165.5 PMOS
M$96 18 20 14 14 PMOS L=1U W=300U AS=420P AD=420P PS=434U PD=434U
* device instance $101 m90 *1 179,165.5 PMOS
M$101 21 21 14 14 PMOS L=1U W=300U AS=360P AD=360P PS=372U PD=372U
* device instance $106 m90 *1 70.5,104.5 PMOS
M$106 3 13 19 19 PMOS L=3U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $111 r0 *1 81.5,104.5 PMOS
M$111 7 8 19 19 PMOS L=3U W=200U AS=240P AD=240P PS=252U PD=252U
* device instance $116 m0 *1 31,123 PMOS
M$116 22 9 19 14 PMOS L=2U W=40U AS=60P AD=60P PS=66U PD=66U
* device instance $118 r180 *1 22,123 PMOS
M$118 24 9 9 14 PMOS L=2U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $123 r0 *1 25,200.5 HRES
R$123 14 1 801500 HRES
* device instance $126 r0 *1 269.75,58 CAP
C$126 18 11 9.49e-13 CAP
* device instance $128 m0 *1 269.25,172.5 CAP
C$128 18 20 9.49e-13 CAP
.ENDS Op8_22_rev2
