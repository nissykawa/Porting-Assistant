* Created by KLayout

* cell Op8_16_rev2
* pin Voutput
* pin Ibias1
* pin In+
* pin In-
* pin Vss
.SUBCKT Op8_16_rev2 7 9 13 17 18
* net 7 Voutput
* net 9 Ibias1
* net 13 In+
* net 17 In-
* net 18 Vss
* device instance $1 r0 *1 219.75,40.2 CAP
C$1 7 5 1.0366e-12 CAP
* device instance $5 r0 *1 55.5,100.5 NMOS
M$5 10 13 12 18 NMOS L=2U W=40U AS=80P AD=80P PS=84U PD=84U
* device instance $6 m90 *1 67.4,100.5 NMOS
M$6 14 17 12 18 NMOS L=2U W=40U AS=80P AD=80P PS=84U PD=84U
* device instance $7 m90 *1 17.1,18.1 NMOS
M$7 3 1 18 18 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $8 r0 *1 28,18.1 NMOS
M$8 2 1 18 18 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $9 r0 *1 113.5,23 NMOS
M$9 5 6 18 18 NMOS L=3U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $10 m90 *1 105,23 NMOS
M$10 6 6 18 18 NMOS L=3U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $11 r0 *1 64.7,35.9 NMOS
M$11 12 1 2 18 NMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $15 m90 *1 57.2,35.9 NMOS
M$15 1 1 3 18 NMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $19 r0 *1 126.3,19.35 NMOS
M$19 7 5 18 18 NMOS L=1U W=25U AS=37.5P AD=37.5P PS=43.5U PD=43.5U
* device instance $21 r0 *1 140.5,127.1 PMOS
M$21 7 9 11 11 PMOS L=5U W=90U AS=120P AD=120P PS=128U PD=128U
* device instance $24 r0 *1 22.6,82.9 PMOS
M$24 1 9 16 11 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $28 r0 *1 121.4,84.7 PMOS
M$28 5 9 10 11 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $32 r0 *1 87.5,84 PMOS
M$32 6 9 14 11 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $36 m90 *1 15,82.9 PMOS
M$36 9 9 15 11 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $40 r0 *1 97.7,127.1 PMOS
M$40 14 9 11 11 PMOS L=5U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $41 r0 *1 24,127 PMOS
M$41 16 9 11 11 PMOS L=5U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $42 m90 *1 13.1,127 PMOS
M$42 15 9 11 11 PMOS L=5U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $43 r0 *1 121,127.1 PMOS
M$43 10 9 11 11 PMOS L=5U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $46 r0 *1 -7.1,31.2 HRES
R$46 18 9 174000 HRES
.ENDS Op8_16_rev2
