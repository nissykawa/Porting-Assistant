* Created by KLayout

* cell TOP
* pin Voutput
* pin Ibias1
* pin Vdd
* pin In+
* pin In-
* pin Vss
.SUBCKT TOP 6 7 9 12 13 16
* net 6 Voutput
* net 7 Ibias1
* net 9 Vdd
* net 12 In+
* net 13 In-
* net 16 Vss
* device instance $1 m90 *1 17.1,18.1 NMOS
M$1 16 1 4 16 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $2 r0 *1 28,18.1 NMOS
M$2 16 1 3 16 NMOS L=5U W=10U AS=20P AD=20P PS=24U PD=24U
* device instance $3 r0 *1 113.5,23 NMOS
M$3 16 5 2 16 NMOS L=3U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $4 m90 *1 105,23 NMOS
M$4 16 5 5 16 NMOS L=3U W=20U AS=40P AD=40P PS=44U PD=44U
* device instance $5 r0 *1 64.7,36 NMOS
M$5 3 1 10 16 NMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $9 m90 *1 57.2,35.9 NMOS
M$9 4 1 1 16 NMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $13 r0 *1 159.2,19.35 NMOS
M$13 16 2 6 16 NMOS L=1U W=25U AS=37.5P AD=37.5P PS=43.5U PD=43.5U
* device instance $15 r0 *1 55.5,100.5 NMOS
M$15 10 12 8 16 NMOS L=2U W=40U AS=80P AD=80P PS=84U PD=84U
* device instance $16 m90 *1 67.4,100.5 NMOS
M$16 10 13 11 16 NMOS L=2U W=40U AS=80P AD=80P PS=84U PD=84U
* device instance $17 r0 *1 140.5,127.1 PMOS
M$17 9 7 6 9 PMOS L=5U W=90U AS=120P AD=120P PS=128U PD=128U
* device instance $20 r0 *1 24,127 PMOS
M$20 9 7 15 9 PMOS L=5U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $21 m90 *1 13.1,127 PMOS
M$21 9 7 14 9 PMOS L=5U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $22 r0 *1 121,127.1 PMOS
M$22 9 7 8 9 PMOS L=5U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $23 r0 *1 97.7,127.1 PMOS
M$23 9 7 11 9 PMOS L=5U W=30U AS=60P AD=60P PS=64U PD=64U
* device instance $24 r0 *1 22.6,82.9 PMOS
M$24 15 7 1 9 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $28 r0 *1 121.4,84.7 PMOS
M$28 8 7 2 9 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $32 r0 *1 87.5,84 PMOS
M$32 11 7 5 9 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $36 m90 *1 15,82.9 PMOS
M$36 14 7 7 9 PMOS L=2U W=100U AS=125P AD=125P PS=135U PD=135U
* device instance $40 r270 *1 136.8,36.6 CAP
C$40 6 2 1.04e-12 CAP
.ENDS TOP
